/*
  CSR ��� ������� � LCD
*/

/* CONTROL REGISTERS */

`define LCD_VER 16'h0_0_0_1

// ������, ������������ �� ���������� ��������� � ILI9341, 
// ����� ������� ���������� �� CPU
`define LCD_DATA_CR      0


// ����������� �������, ������������ �� ���������� ��������� � ILI9341, 
// ����� ������� ���������� �� CPU
`define LCD_CTRL_CR      1
        `define LCD_CTRL_CR_RD      0
        `define LCD_CTRL_CR_WR      1
        `define LCD_CTRL_CR_RS      2

// ���������� ����������
// ���� � ���� �������� ��� ���� ����� 0, �� ������� 
// ���������� �� CPU.
`define LCD_DMA_CR       2
        // ����� ��� ���������� ����������� ���������
        // ����������� ����������� �� LCD
        `define LCD_DMA_CR_REDRAW_STB       0

        // ��������� ����������� (� ������ �������� �������� LCD_FPS_DELAY_CR)
        // ��������� ����������� ����������� �� LCD
        `define LCD_DMA_CR_REDRAW_EN        2

// ������ ����� �����������
`define LCD_DMA_ADDR_CR0 3       
`define LCD_DMA_ADDR_CR1 4

// �������� ����� �����������, � �������������.
// ��������, ������ 25 � ���� ������� ���� 40 FPS.
// ���� �������� �������� ����� 0 
// (��� �����, ���� CPU �� ������� � ������� ������),
// �� ����� ������������ �������� 40 (�� ���� 25 FPS)
`define LCD_FPS_DELAY_CR 5

`define LCD_CR_CNT            6


/* STATUS REGISTERS */

`define LCD_VER_SR 0


`define LCD_DMA_SR 1
        // ��� ����������, ��� ����������� ���������� ������ ������ �� DMA 
        // �� ����������� � ������ �� � LCD.
        // �� ���� ����������� � ILI9341 ������ ��������� FPGA.
        `define LCD_DMA_SR_BUSY 0

`define LCD_SR_CNT 2


/* �������� ������ � LCD-DMA 

  ���� ������ ��������� ���������� ������ �� �����������
  � �������������� DMA � �������� �� �� ILI9341 LCD.

  ����� ������������� ����������� ������� ���������� 
  ���������� ����������� ILI9341 (data, wr, rd, rs).

  ����� ����, ��� ������ ��������� ����������� � ILI9341,
  FPGA ��� CPU, �������������� ��� ������ �������� LCD_DMA_CR.

  �������� 3 ��������:
     * ���������� � CPU
     * ����������� ��������� ����� FPGA
     * ����������� ��������� ����� FPGA (���������� � FPGA)
  
  �� ��������� ���������� ������ CPU.

  ������� ������ (�� ���� 0, ����� 1) � LCD_DMA_CR.LCD_DMA_CR_REDRAW_STB
  �������� � ����, ��� FPGA ���� ��� �������� ������ �� ����������� 
  � ������� �� � LCD.
  �� ������ ���������� ���������� LCD_DMA_SR.LCD_DMA_SR_BUSY ����� ����� 1.

  ������ 1 � LCD_DMA_CR.LCD_DMA_CR_REDRAW_EN �������� � ����, ��� FPGA
  ����� ��������� ���������� ������ �� ����������� � ������ �� � LCD.
  �� �ӣ ����� LCD_DMA_SR.LCD_DMA_SR_BUSY ����� ����� 1.

  ������ ����� ����������� ������ ���� ������� � LCD_DMA_ADDR_CR1/CR0.
  ����� ����� ������ ������ �����, ����� ���������� � CPU.

  �������� �������� FPS � ������� FPGA ����� ������������ ����� 
  � ����������� ������. ��� ����� ����� �������� � ������� LCD_FPS_DELAY_CR 
  �������� (� �������������) ����� ����� ����������� �����. 
  ��������, ������� 25 �� ������� FPS, ������ 40. 
  ���� ������ �� ����������, �� ��������� FPS ����� 25.

*/


